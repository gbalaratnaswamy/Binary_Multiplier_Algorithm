module wallace_multiplier(output [15:0] ans,
input [7:0] m,r
);
wire [7:0] p0,p1,p2,p3,p4,p5,p6,p7;
endmodule


module half_adder (
    output s,cout,
    input a,b
);
    
endmodule


module full_adder (
    output s,cout,
    input a,b,cin
);
    
endmodule